module BullsCows(
    input [15:0] SW,
    input clock,
    input reset,
    input ssl,

    output reg [5:0] d1, d2, d3, d4, d5, d6, d7, d8,
    output reg p1_win,
    output reg p2_win
);
    typedef enum logic [2:0] {S1, S2, T1, T2, RESULT, WIN} state_t;
    state_t state;

    reg [15:0] secret1, secret2;
    integer bulls_int, cows_int;
    reg flag_winner;  // 0: p1, 1: p2

    wire enter_rising;

    edge_detector_s ed (
        .clock(clock),
        .reset(reset),
        .din(ssl),
        .rising(enter_rising)
    );

    // Função para conversão de inteiro para formato 6 bits do display
    function automatic [5:0] to_disp6(input integer value);
        if (value >= 0 && value <= 9)
            to_disp6 = {1'b0, value[3:0], 1'b0};  // enable=0 (ativo), ponto=0
        else
            to_disp6 = 6'h10; // apagado
    endfunction

    // Função de cálculo
    task automatic calc_bulls_cows(
        input [15:0] secret, input [15:0] guess,
        output integer bulls_out, output integer cows_out
    );
        integer i, j;
        reg [3:0] s_digit [3:0], g_digit [3:0];
        bulls_out = 0;
        cows_out = 0;
        for (i = 0; i < 4; i++) begin
            s_digit[i] = secret[i*4 +: 4];
            g_digit[i] = guess[i*4 +: 4];
        end
        for (i = 0; i < 4; i++)
            if (s_digit[i] == g_digit[i]) bulls_out++;
        for (i = 0; i < 4; i++)
            for (j = 0; j < 4; j++)
                if (i != j && s_digit[i] == g_digit[j]) cows_out++;
    endtask

    always_ff @(posedge clock or posedge reset) begin
        if (reset) begin
            state <= S1;
            secret1 <= 0; 
            secret2 <= 0;
            bulls_int <= 0; 
            cows_int <= 0;
            p1_win <= 0; 
            p2_win <= 0;
            flag_winner <= 0;

            d1 <= 6'b111111;  // -
            d2 <= 6'b111111;  // -
            d3 <= 6'b111111;  // -
            d4 <= 6'b111111;  // -
            d5 <= 6'b111111;  // -
            d6 <= 6'b111111;  // -
            d7 <= 6'b111111;  // -
            d8 <= 6'b111111;  // -

        end else begin
            // Limpa pulso após 1 ciclo
            p1_win <= 0;
            p2_win <= 0;

            case (state)
                S1: begin
                    d1 <= 6'hF;  // U
                    d2 <= 6'hD;  // S
                    d3 <= 6'b111111; // -
                    d4 <= 6'h1;  // 1
                    d5 <= 6'hA;  // P
                    d6 <= 6'b111111; // -
                    d7 <= 6'b111111; // -
                    d8 <= 6'b111111; // -
                    if (enter_rising) begin secret1 <= SW; state <= S2; end
                end
                S2: begin
                    d1 <= 6'hF;  // U
                    d2 <= 6'hD;  // S
                    d3 <= 6'b111111; // -
                    d4 <= 6'h2;  // 2
                    d5 <= 6'hA;  // P
                    d6 <= 6'b111111; // -
                    d7 <= 6'b111111; // -
                    d8 <= 6'b111111; // -
                    if (enter_rising) begin secret2 <= SW; state <= T1; end
                end
                T1: begin
                    d1 <= 6'h6;  // G (6)
                    d2 <= 6'b111111; // -
                    d3 <= 6'h1;  // 1
                    d4 <= 6'hA;  // P
                    d5 <= 6'b111111; // -
                    d6 <= 6'b111111; // -
                    d7 <= 6'b111111; // -
                    d8 <= 6'b111111; // -
                    if (enter_rising) begin
                        calc_bulls_cows(secret2, SW, bulls_int, cows_int);
                        if (bulls_int == 4) begin flag_winner <= 0; state <= WIN; end
                        else state <= RESULT;
                    end
                end
                T2: begin
                    d1 <= 6'h6;  // G (6)
                    d2 <= 6'b111111; // -
                    d3 <= 6'h2;  // 1
                    d4 <= 6'hA;  // P
                    d5 <= 6'b111111; // -
                    d6 <= 6'b111111; // -
                    d7 <= 6'b111111; // -
                    d8 <= 6'b111111; // -
                    if (enter_rising) begin
                        calc_bulls_cows(secret1, SW, bulls_int, cows_int);
                        if (bulls_int == 4) begin flag_winner <= 1; state <= WIN; end
                        else state <= RESULT;
                    end
                end
                RESULT: begin
                    d1 <= to_disp6(bulls_int); // número de touros
                    d2 <= 6'hB;                // letra "b"
                    d3 <= 6'h10;               // -
                    d4 <= to_disp6(cows_int);  // número de vacas
                    d5 <= 6'hC;                // letra "c"
                    d6 <= 6'b111111;           // -
                    d7 <= 6'b111111;           // -
                    d8 <= 6'b111111;           // -
                    if (enter_rising) begin
                        bulls_int <= 0;
                        cows_int <= 0;
                        state <= (flag_winner == 0) ? T2 : T1;
                    end
                end
                WIN: begin
                    d1 <= 6'hE;  // E  
                    d2 <= 6'b111111; // -
                    d3 <= 6'hB;  // B
                    d4 <= 6'b111111; // -
                    d5 <= 6'b111111; // -
                    d6 <= 6'b111111; // -
                    d7 <= 6'b111111; // -
                    d8 <= 6'b111111; // -
                    if (flag_winner == 0) p1_win <= 1;
                    else p2_win <= 1;
                    if (enter_rising) state <= S1;
                end
            endcase
        end
    end
endmodule
