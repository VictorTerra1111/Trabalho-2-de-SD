module switch(
    input logic sw[15:0],
    output logic out[15:0]
);

assign out = sw;

endmodule
