module switch(
input logic sw,
output logic out

);

assign out = sw;

endmodule
